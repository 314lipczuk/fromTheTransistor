
module test 
// port list
	(
	in_1,
	in_2,
	out_1,
	carry
	);
// port & wire definition
	input	in_1;
	input	in_2;
	output 	out_1;
	output 	carry;

// Implementation & assigning wires 
//
//
endmodule


// assign s are continuous - they work simultaneously, have no memory, and
// rely only on inputs at a given time (direct combinatorial logic)


