module blink_led

endmodule
